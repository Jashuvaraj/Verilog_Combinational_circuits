module Full_adder_tb;
reg a,b,c;
wire s,cin;
Full_adder dut(a,b,c,s,cin);
initial begin
#10 a=0;b=0;c=0;
#10 a=0;b=0;c=1;
#10 a=0;b=1;c=0;
#10 a=0;b=1;c=1;
#10 a=1;b=0;c=0;
#10 a=1;b=0;c=1;
#10 a=1;b=1;c=0;
#10 a=1;b=1;c=1;
end 
endmodule
